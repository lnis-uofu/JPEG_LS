`timescale 1ns/1ns
`include "Parameterize_JPEGLS.v"
/* 
======================================================================================================================================================================================================
	AUTHOR: GRANT BROWN (LNIS)
	DATE: 4/18/2020
	DESCRIPTION: The K value is a Golomb coding parameter. Value is calcualted within this module. The max value for k is 14 due to the max value of A being 8191. Priority based architecture
		     used in this module due to the nature of sequential operation.
======================================================================================================================================================================================================
*/
module k_calculation_unrolled #(parameter N_length = `N_length, A_length = `A_length, mode_length = `mode_length, temp_length = `temp_length, k_length = `k_length)
		     	       (input [N_length - 1 : 0] N, input [A_length - 1 : 0] A, input [mode_length - 1 : 0] mode, input RIType, 
		       		input [temp_length  - 1 : 0] temp, input [k_length - 1: 0] k_inc, output reg [k_length - 1:0] k);

/* 
======================================================================================================================================================================================================
	WIRE DECLARATION
======================================================================================================================================================================================================
*/

	reg [k_length - 1:0] k_index;
	wire [k_length - 1:0] k_RGM;
	wire [k_length - 1:0] k_RIM;

/* 
======================================================================================================================================================================================================
	REG DECLARATION
======================================================================================================================================================================================================
*/
	defparam Regular_Mode_K.Iteration_Count = 14;
	K_Determination Regular_Mode_K (.A(A), .N(N), .k_index(k_inc), .k(k_RGM));

/* 
======================================================================================================================================================================================================
	MODULE INSTANTIATION
======================================================================================================================================================================================================
*/

	defparam Run_Interrupt_K.A_length = temp_length;
	K_Determination Run_Interrupt_K (.A(temp), .N(N), .k_index(k_inc), .k(k_RIM));

/* 
======================================================================================================================================================================================================
	COMBINATIONAL LOGIC
======================================================================================================================================================================================================
*/

	always @ (N or A or mode or RIType or temp or k_RIM or k_RGM) begin
		k_index = k_inc;
		k = k_inc;
		if (mode == 0) begin
			k = k_RGM;
		end
		// run interruption coding
		else if (mode == 2) begin
			k = k_RIM;
		end
		else k = 0;
	end


endmodule