`timescale 1ns/1ns
`include "Parameterize_JPEGLS.v"
/* 
======================================================================================================================================================================================================
	AUTHOR: GRANT BROWN (LNIS)
	DATE: 4/18/2020
	DESCRIPTION: Updates N value and determiens if N needs to be reset based on variable threshold value. Hides the reset from stalling the pipeline.
======================================================================================================================================================================================================
*/
module NUpdate #(parameter N_length = `N_length)
		(input [N_length - 1:0] N, output reg resetFlag, output reg [N_length - 1:0] N_New);

/* 
======================================================================================================================================================================================================
	GENERALIZED PARAMETER DECLARATIONS
======================================================================================================================================================================================================
*/
	localparam [N_length - 1:0] threshold = 64;

/* 
======================================================================================================================================================================================================
	COMBINATIONAL LOGIC
======================================================================================================================================================================================================
*/

	always @ (N) begin
		if (N == threshold) begin
			N_New = (N >> 1) + 1;
			resetFlag = 1;
		end
		else begin
			N_New = N + 1;
			resetFlag = 0;
		end
	end
endmodule
