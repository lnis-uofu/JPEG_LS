`timescale 1ns/1ns
`include "Parameterize_JPEGLS.v"

/* 
======================================================================================================================================================================================================
	AUTHOR: GRANT BROWN (LNIS)
	DATE: 7/7/2020
	DESCRIPTION: Internal calculation module for the Golomb k value. The iteration count is fixed therefore the for loop is synthesizable. Follows the standard set forth by the ITU T.87
======================================================================================================================================================================================================
*/

module K_Determination (A, N, k_index, k);

/* 
======================================================================================================================================================================================================
	GENERALIZED PARAMETER DECLARATIONS
======================================================================================================================================================================================================
*/

	parameter A_length = `A_length;
	parameter Iteration_Count = 15;
	localparam N_length = `N_length;
	localparam k_length = `k_length;

/* 
======================================================================================================================================================================================================
	REG DECLARATION
======================================================================================================================================================================================================
*/

	integer k_inc, temp;

/* 
======================================================================================================================================================================================================
	I/O DECLARATION
======================================================================================================================================================================================================
*/

	input [A_length - 1:0] A;
	input [N_length - 1:0] N;
	input [k_length - 1:0] k_index;
	output reg [k_length - 1:0] k;

/* 
======================================================================================================================================================================================================
	COMBINATIONAL LOGIC
======================================================================================================================================================================================================
*/


	always @ (A or N or k_index) begin
		k = k_index;
		for(k_inc  = 0; k_inc < Iteration_Count; k_inc = k_inc + 1) begin
			temp = N << k_inc;
			if (temp < A) k = k + 1;
			else k = k;
		end
	end

endmodule
